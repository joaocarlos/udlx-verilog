// +----------------------------------------------------------------------------
// GNU General Public License
// -----------------------------------------------------------------------------
// This file is part of uDLX (micro-DeLuX) soft IP-core.
//
// uDLX is free soft IP-core: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// uDLX soft core is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with uDLX. If not, see <http://www.gnu.org/licenses/>.
// +----------------------------------------------------------------------------
// PROJECT: uDLX core Processor
// ------------------------------------------------------------------------------
// FILE NAME        : config.vh
// AUTHOR(s)        : joaocarlos
// MANTAINER        : joaocarlos
// AUTHOR'S E-MAIL  : joaocarlos@ieee.org
// -----------------------------------------------------------------------------
// KEYWORDS: parameters, config, dlx
// -----------------------------------------------------------------------------
// PURPOSE: IP core header configuration file
// -----------------------------------------------------------------------------


// -------------------------------------------------------------
// Main configuration
// -------------------------------------------------------------
`define CORE_WIDTH 32

// -------------------------------------------------------------
// Opcodes
// -------------------------------------------------------------
// Arithmetical Logic Unit
`define ADD
`define SUB
`define AND
`define OR
`define MULT
`define DIV
`define CMP
`define NOT

// -------------------------------------------------------------
// Flags
// -------------------------------------------------------------