clk_40_inst : clk_40 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
